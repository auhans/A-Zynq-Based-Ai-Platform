`timescale 1ns / 1ps


module vmx_execute_processor(
    input wire [31:0] test,
    output reg [31:0] test2
    );
endmodule
